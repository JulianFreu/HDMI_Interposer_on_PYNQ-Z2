attribute ram_style : string;
attribute ram_style of myram : signal is "ultra";
